/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 919;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_656e6f64,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d79726f_6d656d20,
        64'h6e69616d_206f7420,
        64'h00000020_6874676e,
        64'h656c2068_74697720,
        64'h00000020_6d6f7266,
        64'h20676e69_79706f43,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00322d74_6c756166,
        64'h65642d69_72742c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_6972742c,
        64'h786e6c78_006c6175,
        64'h642d7369_2c786e6c,
        64'h7800746e_65736572,
        64'h702d7470_75727265,
        64'h746e692c_786e6c78,
        64'h00687464_69772d32,
        64'h6f697067_2c786e6c,
        64'h78006874_6469772d,
        64'h6f697067_2c786e6c,
        64'h7800322d_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800746c,
        64'h75616665_642d7475,
        64'h6f642c78_6e6c7800,
        64'h322d7374_75706e69,
        64'h2d6c6c61_2c786e6c,
        64'h78007374_75706e69,
        64'h2d6c6c61_2c786e6c,
        64'h78007265_6c6c6f72,
        64'h746e6f63_2d6f6970,
        64'h6700736c_6c65632d,
        64'h6f697067_23007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_ad020000,
        64'h04000000_03000000,
        64'hffffffff_9c020000,
        64'h04000000_03000000,
        64'h01000000_8f020000,
        64'h04000000_03000000,
        64'h00000000_78020000,
        64'h04000000_03000000,
        64'h08000000_67020000,
        64'h04000000_03000000,
        64'h08000000_57020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_1f020000,
        64'h04000000_03000000,
        64'h00000000_0f020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_ff010000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'hf3010000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h03000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h30080000_c0020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h68080000_38000000,
        64'h280b0000_edfe0dd0,
        64'h33323130_2f2e2d2c,
        64'h2b2a2928_27262524,
        64'h23222120_1f1e1d1c,
        64'h1b1affff_ffffffff,
        64'h19181716_15141312,
        64'h11100f0e_0d0c0b0a,
        64'h09080706_05040302,
        64'h0100ffff_fffeffff,
        64'hff3d3c3b_3a393837,
        64'h3635343f_ffffff3e,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'ha0018402_17458593,
        64'h00000597_01f41413,
        64'h0010041b_cb0ff0ef,
        64'hd0050513_00001517,
        64'hff2491e3_87a6cc2f,
        64'hf0efd0a5_05130000,
        64'h1517e799_0084f7b3,
        64'hc39897ce_00478493,
        64'h43986200_0937147d,
        64'h1f0009b7_610007b7,
        64'h00080437_cf0ff0ef,
        64'hd2050513_00001517,
        64'hd94ff0ef_01000537,
        64'hd04ff0ef_d2450513,
        64'h00001517_da8ff0ef,
        64'h61000537_d18ff0ef,
        64'hd2850513_00001517,
        64'hd24ff0ef_d2450513,
        64'h00001517_cecff0ef,
        64'hec26e44e_e84af022,
        64'hf4060805_05132005,
        64'h85937179_02faf537,
        64'h65f1bdf5_00aa8023,
        64'h8d5d03f5_7513000a,
        64'hc783e9bf_f0ef001a,
        64'h84930014_8a130004,
        64'hc503bf15_00f90223,
        64'h408a853b_000ac783,
        64'h00f92023_478d00f4,
        64'h9c630169_87b300aa,
        64'h00a300fa_00230065,
        64'h151b8fd9_8bbd4025,
        64'h579b000a_4703edff,
        64'hf0ef001a_0a93001a,
        64'h8493000a_c503b7c5,
        64'h8aaa8a32_bfbd00f9,
        64'h0223408a_053b000a,
        64'h478300f9_20234789,
        64'h00fa9f63_016987b3,
        64'h00a480a3_00f48023,
        64'h0045151b_8fd98b8d,
        64'h4045579b_0004c703,
        64'hf29ff0ef_00148a13,
        64'h001b8a93_000bc503,
        64'hb7f58baa_84b2bf75,
        64'h00f92023_478500fb,
        64'h99630169_87b300a4,
        64'h80230025_151bf57f,
        64'hf0ef001a_0b93000a,
        64'h45038082_61616ba2,
        64'h6b426ae2_7a0279a2,
        64'h794274e2_640660a6,
        64'h00f90223_4084853b,
        64'h0004c783_00092023,
        64'h02fa1563_016987b3,
        64'h8a2a84b2_a8c184ce,
        64'h8ab202e7_93634501,
        64'h470d0ae7_89634709,
        64'hcb9906e7_88638936,
        64'h84328b2e_89aa4705,
        64'he45eec56_f052fc26,
        64'he486e85a_f44ef84a,
        64'h429c00f6_0023e0a2,
        64'h715d0046_c7838082,
        64'h00050223_00052023,
        64'h8082557d_80820007,
        64'hc50397aa_33478793,
        64'h00000797_00a7ea63,
        64'h04f00793_0ff57513,
        64'hfd55051b_b38decaf,
        64'hf0ef1fa5_05130000,
        64'h1517bbd9_f5c50513,
        64'h00001517_f78ff0ef,
        64'h8526ee6f_f0ef0565,
        64'h05130000_1517ef2f,
        64'hf0ef04a5_05130000,
        64'h1517bbfd_f8450513,
        64'h00001517_fa0ff0ef,
        64'h8526f0ef_f0ef07e5,
        64'h05130000_1517f1af,
        64'hf0ef0725_05130000,
        64'h1517c929_84aac3df,
        64'hf0ef8556_865e020b,
        64'h2583f36f_f0ef24e5,
        64'h05130000_1517f384,
        64'h9de30809_0913080a,
        64'h0993f4ef_f0ef2485,
        64'hfd850513_00001517,
        64'hff3a1be3_83bff0ef,
        64'h0a05000a_4503f6af,
        64'hf0ef2725_05130000,
        64'h151780ff_f0ef0109,
        64'h3503f7ef_f0ef2765,
        64'h05130000_1517823f,
        64'hf0ef0089_3503f92f,
        64'hf0ef27a5_05130000,
        64'h1517837f_f0effb89,
        64'h8a130009_3503faaf,
        64'hf0ef2825_05130000,
        64'h1517ff2a_1be3895f,
        64'hf0ef0a05_000a4503,
        64'hf9098a13_fc8ff0ef,
        64'h28050513_00001517,
        64'hff9a19e3_8b3ff0ef,
        64'h0a050007_c503014d,
        64'h07b34a01_fe8ff0ef,
        64'hf8098d13_28450513,
        64'h00001517_8d3ff0ef,
        64'h0ff4f513_801ff0ef,
        64'h28050513_00001517,
        64'h4c114cc1_10051b63,
        64'h02010913_08010993,
        64'h84aa8b0a_d33ff0ef,
        64'h850a4605_71010489,
        64'h258382ff_f0ef0b65,
        64'h05130000_1517893f,
        64'hf0ef4556_841ff0ef,
        64'h2a050513_00001517,
        64'h8a5ff0ef_4546853f,
        64'hf0ef2925_05130000,
        64'h15178f7f_f0ef6526,
        64'h865ff0ef_28450513,
        64'h00001517_909ff0ef,
        64'h7502877f_f0ef2865,
        64'h05130000_151791bf,
        64'hf0ef6562_889ff0ef,
        64'h28050513_00001517,
        64'h8edff0ef_455289bf,
        64'hf0ef2825_05130000,
        64'h15178fff_f0ef4542,
        64'h8adff0ef_28450513,
        64'h00001517_911ff0ef,
        64'h45328bff_f0ef2865,
        64'h05130000_1517923f,
        64'hf0ef4522_8d1ff0ef,
        64'h28850513_00001517,
        64'h975ff0ef_65028e3f,
        64'hf0ef28a5_05130000,
        64'h15178eff_f0ef2765,
        64'h05130000_1517bf51,
        64'h54f98fff_f0ef1865,
        64'h05130000_15179a3f,
        64'hf0ef8526_911ff0ef,
        64'h28050513_00001517,
        64'h91dff0ef_27450513,
        64'h00001517_c90584aa,
        64'h890ae41f_f0ef850a,
        64'h45854605_710193bf,
        64'hf0ef27a5_05130000,
        64'h15178082_61256d02,
        64'h6ca26c42_6be27b02,
        64'h7aa27a42_79e26906,
        64'h64a66446_852660e6,
        64'hfa040113_54fd96bf,
        64'hf0ef2825_05130000,
        64'h1517c90d_defff0ef,
        64'h8bae8aaa_1080e06a,
        64'he466e862_f05af852,
        64'hfc4ee0ca_e4a6ec86,
        64'hec5ef456_e8a2711d,
        64'hb7655479_80826169,
        64'h6baa6b4a_6aea7a0a,
        64'h79aa794a_74ea640e,
        64'h60ae8522_547d9bbf,
        64'hf0ef2b25_05130000,
        64'h1517c5df_f0efc61f,
        64'hf0efc65f_f0efc69f,
        64'hf0efc6df_f0efc71f,
        64'hf0efc75f_f0efc79f,
        64'hf0efa805_c7fff0ef,
        64'hc8bff0ef_45314581,
        64'h46054401_f93046e3,
        64'h20048493_19fda03f,
        64'hf0ef24a5_05130000,
        64'h1517e799_0369e7b3,
        64'h06891c63_90412901,
        64'h14428c49_cb7ff0ef,
        64'h90410305_14130085,
        64'h151bcc5f_f0effc94,
        64'h1ae30404_0413ff7a,
        64'h17e3892a_f15ff0ef,
        64'h0a05854a_0007c583,
        64'h014407b3_04000b93,
        64'h4a01c69f_f0ef850a,
        64'h04000593_86224901,
        64'hff551ee3_cffff0ef,
        64'he0048413_3e800b13,
        64'h0fe00a93_e9512004,
        64'h8493d1df_f0ef4549,
        64'h85a20ff6_76130016,
        64'h66130015_161bf4df,
        64'hf0ef0ff4_7593f55f,
        64'hf0ef0ff5_f5930084,
        64'h559bf61f_f0ef0ff5,
        64'hf5930104_559bf6df,
        64'hf0ef4501_0184559b,
        64'hfee79be3_078500c6,
        64'h802300f1_06b30800,
        64'h0713567d_47810209,
        64'hd993842e_84aae55e,
        64'he95aed56_f152f94a,
        64'he586fd26_e1a20206,
        64'h1993f54e_71558082,
        64'h91411542_8d3d8ff9,
        64'h0057979b_17016709,
        64'h0107d79b_0105179b,
        64'h4105551b_0105151b,
        64'h8d2d00c5_95138da9,
        64'h893d0045_d51b8da9,
        64'h91411542_8d5d0522,
        64'h0085579b_808207f5,
        64'h75138d2d_00451593,
        64'h8d2d8d3d_0045d51b,
        64'h0075d79b_8de98082,
        64'h0141853e_640260a2,
        64'h57f5e111_4781f89f,
        64'hf0efc511_57f9efbf,
        64'hf0efc911_57fdeb7f,
        64'hf0effc6d_e07ff0ef,
        64'h347d4429_b79ff0ef,
        64'h45850513_00001517,
        64'hc89ff0ef_e022e406,
        64'h11418082_61050015,
        64'h351364a2_644260e2,
        64'h0004051b_fc940ce3,
        64'he3bff0ef_eb3ff0ef,
        64'h48050513_00001517,
        64'h85aa842a_e57ff0ef,
        64'h02900513_400005b7,
        64'h07700613_fbdff0ef,
        64'h4485e822_ec06e426,
        64'h11018082_01410015,
        64'h3513157d_640260a2,
        64'h0004051b_ef3ff0ef,
        64'h4ba50513_85a20000,
        64'h1517e8df_f0ef842a,
        64'he9bff0ef_e022e406,
        64'h03700513_45810650,
        64'h06131141_80826105,
        64'h690264a2_644260e2,
        64'h00153513_f5650513,
        64'h0004051b_01249863,
        64'h88bd00f9_1b634501,
        64'h4785ecdf_f0efed1f,
        64'hf0ef842a_ed7ff0ef,
        64'h84aaeddf_f0efee1f,
        64'hf0efee5f_f0ef892a,
        64'hef3ff0ef_e04ae426,
        64'he822ec06_45211aa0,
        64'h05930870_06131101,
        64'hbfcd4501_80826105,
        64'h690264a2_644260e2,
        64'h4505f89f_f0ef4585,
        64'h54850513_00001517,
        64'hfe9915e3_c00df29f,
        64'hf0ef892a_347df39f,
        64'hf0ef4501_45810950,
        64'h06134485_71040413,
        64'he04aec06_e4266409,
        64'he8221101_cb9ff06f,
        64'h61055425_05130000,
        64'h151760e2_6442da5f,
        64'hf0ef852e_65a2cd3f,
        64'hf0ef58a5_05130000,
        64'h1517cdff_f0ef8522,
        64'hce5ff0ef_e42eec06,
        64'h59050513_00001517,
        64'h842ae822_11018082,
        64'h614564e2_740270a2,
        64'hf47d147d_0007d463,
        64'h4187d79b_0185179b,
        64'hfabff0ef_eb5ff0ef,
        64'h85320640_04136622,
        64'hec1ff0ef_0ff47513,
        64'hec9ff0ef_0ff57513,
        64'h0084551b_ed5ff0ef,
        64'h0ff57513_0104551b,
        64'hee1ff0ef_0184551b,
        64'hee9ff0ef_0404e513,
        64'hfebff0ef_84aa842e,
        64'hec26f022_e432f406,
        64'h7179f03f_f06f0ff0,
        64'h05138082_557db7d9,
        64'h00d70023_078500f6,
        64'h073306c8_2683ff69,
        64'h8b055178_b77dd6b8,
        64'h07850007_470300f5,
        64'h07338082_4501d3b8,
        64'h4719dbb8_577d2000,
        64'h07b702b6_e1630007,
        64'h869b2000_08372000,
        64'h0537fff5_8b85537c,
        64'h20000737_d3b82000,
        64'h07b71060_0713fff5,
        64'h37fd0001_03200793,
        64'h04b76163_0007871b,
        64'h47812000_06b7dbb8,
        64'h57792000_07b706b7,
        64'hee631000_07938082,
        64'h610564a2_d3b84719,
        64'hdbb86442_60e20ff4,
        64'h7513577d_200007b7,
        64'he0dff0ef_69450513,
        64'h00001517_eb1ff0ef,
        64'h91011502_4088e23f,
        64'hf0ef6b25_05130000,
        64'h1517e395_8b852401,
        64'h53fc57e0_ff658b05,
        64'h06478493_53f8d3b8,
        64'h10600713_200007b7,
        64'hfff537fd_00010640,
        64'h0793d7a8_dbb85779,
        64'he426e822_ec062000,
        64'h07b71101_e69ff06f,
        64'h61056e25_05130000,
        64'h151764a2_60e26442,
        64'hd03c4799_e81ff0ef,
        64'h70850513_00001517,
        64'hf25ff0ef_91010204,
        64'h95132481_e99ff0ef,
        64'h70050513_00001517,
        64'h5064d03c_16600793,
        64'headff0ef_73450513,
        64'h00001517_f51ff0ef,
        64'h91010204_95132481,
        64'hec5ff0ef_72c50513,
        64'h00001517_5064d03c,
        64'h10400793_20000437,
        64'hfff537fd_000147a9,
        64'hc3b84729_200007b7,
        64'heedff0ef_e426e822,
        64'hec0674c5_05131101,
        64'h00001517_80822501,
        64'h41088082_c10c8082,
        64'h610560e2_eb9ff0ef,
        64'h00914503_ec1ff0ef,
        64'h00814503_f55ff0ef,
        64'hec06002c_11018082,
        64'h61456942_64e27402,
        64'h70a2fe94_10e3ee3f,
        64'hf0ef0091_4503eebf,
        64'hf0ef3461_00814503,
        64'hf81ff0ef_0ff57513,
        64'h002c0089_553354e1,
        64'h03800413_892af406,
        64'he84aec26_f0227179,
        64'h80826145_694264e2,
        64'h740270a2_fe9410e3,
        64'hf25ff0ef_00914503,
        64'hf2dff0ef_34610081,
        64'h4503fc3f_f0ef0ff5,
        64'h7513002c_0089553b,
        64'h54e14461_892af406,
        64'he84aec26_f0227179,
        64'h808200f5_80230007,
        64'hc78300e5_80a397aa,
        64'h81110007_4703973e,
        64'h00f57713_b4c78793,
        64'h00001797_f79ff06f,
        64'h80820007_4503dfed,
        64'h8b850147_47831000,
        64'h0737b7f5_0405f93f,
        64'hf0ef8082_01416402,
        64'h60a2e509_00044503,
        64'h842ae406_e0221141,
        64'h808200e7_88230200,
        64'h071300e7_8423fc70,
        64'h071300e7_8623470d,
        64'h00a78223_0ff57513,
        64'h00e78023_0085551b,
        64'h0ff57713_00e78623,
        64'hf8000713_00078223,
        64'h100007b7_02b5553b,
        64'h0045959b_808200a7,
        64'h0023dfe5_0207f793,
        64'h01474783_10000737,
        64'h80828905_0147c503,
        64'h100007b7_80820205,
        64'h75130147_c5031000,
        64'h07b78082_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_dd458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h41b000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
